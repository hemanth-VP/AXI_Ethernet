module readme
endmodule
