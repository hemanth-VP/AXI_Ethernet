module top;
endmodule 
